----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:46:02 08/01/2008 
-- Design Name: 
-- Module Name:    Ram - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
--------------------------------------------------------------------------------------------
-- Dual-Port Block RAM with Different Clocks
-- XST User Guide - RAMs and ROMs HDL Coding Techniques
--------------------------------------------------------------------------------------------
library ieee; use ieee.std_logic_1164.all; use ieee.std_logic_unsigned.all;

entity dpram_t2 is
	generic ( BUS_WIDTH  : integer range 1 to   16 :=   16;		--    8
			    ADDR_WIDTH : integer range 1 to   12 :=   11;		--   12
			    RAM_DEPTH	: integer range 1 to 4096 := 1600); 	-- 3200
	port (clka : in  std_logic;
			clkb : in  std_logic;
			wea  : in  std_logic;
			addra: in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			addrb: in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			dia  : in  std_logic_vector(BUS_WIDTH-1 downto 0);
			doa  : out std_logic_vector(BUS_WIDTH-1 downto 0);
			dob  : out std_logic_vector(BUS_WIDTH-1 downto 0));
end dpram_t2;

architecture syn of dpram_t2 is
	type ram_type is array (RAM_DEPTH-1 downto 0) of std_logic_vector (BUS_WIDTH-1 downto 0);
	signal RAM : ram_type:=
	(
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",


		x"0100",x"0302",x"0504",x"0706",x"0908",x"0b0a",x"0d0c",x"0f0e",x"1110",x"1312",
		x"1514",x"1716",x"1918",x"1b1a",x"1d1c",x"1f1e",x"2120",x"2322",x"2524",x"2726",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",

		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020"

	);
	
	signal read_addra : std_logic_vector(ADDR_WIDTH-1 downto 0);
	signal read_addrb : std_logic_vector(ADDR_WIDTH-1 downto 0);
	begin
		process (clka)	begin
			if (rising_edge(clka)) then
				if (wea = '1') then
					RAM(conv_integer(addra)) <= dia;
				end if;
				read_addra <= addra;
			end if;
		end process;

		process (clkb)	begin
			if (rising_edge(clkb)) then
				read_addrb <= addrb;
			end if;
		end process;
		
		doa <= RAM(conv_integer(read_addra));
		dob <= RAM(conv_integer(read_addrb));
end syn;


------------------------------------------------------------------------------------------
--											End of file
--------------------------------------------------------------------------------------------
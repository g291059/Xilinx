----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:46:02 08/01/2008 
-- Design Name: 
-- Module Name:    Ram - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
--------------------------------------------------------------------------------------------
-- Dual-Port Block RAM with Different Clocks
-- XST User Guide - RAMs and ROMs HDL Coding Techniques
--------------------------------------------------------------------------------------------
library ieee; use ieee.std_logic_1164.all; use ieee.std_logic_unsigned.all;

entity dpram_t2 is
	generic ( BUS_WIDTH  : integer range 1 to   16 :=   16;		--    8
			    ADDR_WIDTH : integer range 1 to   12 :=   11;		--   12
			    RAM_DEPTH	: integer range 1 to 4096 := 1600); 	-- 3200
	port (clka : in  std_logic;
			clkb : in  std_logic;
			wea  : in  std_logic;
			addra: in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			addrb: in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			dia  : in  std_logic_vector(BUS_WIDTH-1 downto 0);
			doa  : out std_logic_vector(BUS_WIDTH-1 downto 0);
			dob  : out std_logic_vector(BUS_WIDTH-1 downto 0));
end dpram_t2;

architecture syn of dpram_t2 is
	type ram_type is array (RAM_DEPTH-1 downto 0) of std_logic_vector (BUS_WIDTH-1 downto 0);
	signal RAM : ram_type:=
	(
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
	
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",

		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938"
	
	);
	
	signal read_addra : std_logic_vector(ADDR_WIDTH-1 downto 0);
	signal read_addrb : std_logic_vector(ADDR_WIDTH-1 downto 0);
	begin
		process (clka)	begin
			if (rising_edge(clka)) then
				if (wea = '1') then
					RAM(conv_integer(addra)) <= dia;
				end if;
				read_addra <= addra;
			end if;
		end process;

		process (clkb)	begin
			if (rising_edge(clkb)) then
				read_addrb <= addrb;
			end if;
		end process;
		
		doa <= RAM(conv_integer(read_addra));
		dob <= RAM(conv_integer(read_addrb));
end syn;

--------------------------------------------------------------------------------------------
-- Dual-Port RAM with One Enable Controlling Both Ports
-- XST User Guide - RAMs and ROMs HDL Coding Techniques
--------------------------------------------------------------------------------------------
--library IEEE;use IEEE.STD_LOGIC_1164.ALL;use IEEE.STD_LOGIC_ARITH.ALL;use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
--entity dpram_t1 is
--	 generic ( BUS_WIDTH  : integer range 1 to   16 :=   16;		--    8
--				  ADDR_WIDTH : integer range 1 to   12 :=   11;		--   12
--				  RAM_DEPTH	 : integer range 1 to 4096 := 1600); 	-- 3200
--    port (  ck    : in  std_logic;
--				en		: in  std_logic;
--				we   	: in  std_logic;
--				addra : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
--				addrb : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
--				di    : in  std_logic_vector(BUS_WIDTH-1 downto 0);
--				doa   : out std_logic_vector(BUS_WIDTH-1 downto 0);
--				dob   : out std_logic_vector(BUS_WIDTH-1 downto 0));
--end dpram_t1;
--
--configuration dpram1 of dpram_t1 is
--	for Width16
--	end for;
--end configuration dpram1;
--
--architecture Behavioral of dpram_t1 is
--	type ram_type is array (0 to RAM_DEPTH-1) of std_logic_vector (BUS_WIDTH-1 downto 0);
--	signal vga_ram : ram_type :=
--	(
--		x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",
--		x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",
--		x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",
--		x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",
--
--
--		x"00",x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"0a",x"0b",x"0c",x"0d",x"0e",x"0f",x"10",x"11",x"12",x"13",
--		x"14",x"15",x"16",x"17",x"18",x"19",x"1a",x"1b",x"1c",x"1d",x"1e",x"1f",x"20",x"21",x"22",x"23",x"24",x"25",x"26",x"27",
--		x"28",x"29",x"2a",x"2b",x"2c",x"2d",x"2e",x"2f",x"30",x"31",x"32",x"33",x"34",x"35",x"36",x"37",x"38",x"39",x"3a",x"3b",
--		x"3c",x"3d",x"3e",x"3f",x"40",x"41",x"42",x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4a",x"4b",x"4c",x"4d",x"4e",x"4f",
--
--		x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57",x"58",x"59",x"5a",x"5b",x"5c",x"5d",x"5e",x"5f",x"60",x"61",x"62",x"63",
--		x"64",x"65",x"66",x"67",x"68",x"69",x"6a",x"6b",x"6c",x"6d",x"6e",x"6f",x"70",x"71",x"72",x"73",x"74",x"75",x"76",x"77",
--		x"78",x"79",x"7a",x"7b",x"7c",x"7d",x"7e",x"7f",x"80",x"81",x"82",x"83",x"84",x"85",x"86",x"87",x"88",x"89",x"8a",x"8b",
--		x"8c",x"8d",x"8e",x"8f",x"90",x"91",x"92",x"93",x"94",x"95",x"96",x"97",x"98",x"99",x"9a",x"9b",x"9c",x"9d",x"9e",x"9f",
--
--		x"a0",x"a1",x"a2",x"a3",x"a4",x"a5",x"a6",x"a7",x"a8",x"a9",x"aa",x"ab",x"ac",x"ad",x"ae",x"af",x"b0",x"b1",x"b2",x"b3",
--		x"b4",x"b5",x"b6",x"b7",x"b8",x"b9",x"ba",x"bb",x"bc",x"bd",x"be",x"bf",x"c0",x"c1",x"c2",x"c3",x"c4",x"c5",x"c6",x"c7",
--		x"c8",x"c9",x"ca",x"cb",x"cc",x"cd",x"ce",x"cf",x"d0",x"d1",x"d2",x"d3",x"d4",x"d5",x"d6",x"d7",x"d8",x"d9",x"da",x"db",
--		x"dc",x"dd",x"de",x"df",x"e0",x"e1",x"e2",x"e3",x"e4",x"e5",x"e6",x"e7",x"e8",x"e9",x"ea",x"eb",x"ec",x"ed",x"ee",x"ef",
--
--		x"f0",x"f1",x"f2",x"f3",x"f4",x"f5",x"f6",x"f7",x"f8",x"f9",x"fa",x"fb",x"fc",x"fd",x"fe",x"ff",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
--		x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20"	
--
--	);
--	signal read_addra : std_logic_vector(ADDR_WIDTH-1 downto 0);
--	signal read_addrb : std_logic_vector(ADDR_WIDTH-1 downto 0);
--begin
--	process (ck)
--	begin
--		if (rising_edge(ck)) then
--			if (en = '1') then
--				if (we = '1') then
--					vga_ram(conv_integer(addra)) <= di;
--				end if;
--				read_addra <= addra;
--				read_addrb <= addrb;
--			end if;
--		end if;
--	end process;
--	doa <= vga_ram(conv_integer(read_addra));
--	dob <= vga_ram(conv_integer(read_addrb));
--end Behavioral;
--------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------
--
--architecture Width16 of dpram_t1 is
--	type ram_type is array (0 to RAM_DEPTH-1) of std_logic_vector (BUS_WIDTH-1 downto 0);
--	signal vga_ram : ram_type :=
--	(
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--
--
--		x"0100",x"0302",x"0504",x"0706",x"0908",x"0b0a",x"0d0c",x"0f0e",x"1110",x"1312",
--		x"1514",x"1716",x"1918",x"1b1a",x"1d1c",x"1f1e",x"2120",x"2322",x"2524",x"2726",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--		x"3130",x"3332",x"3534",x"3736",x"3938",x"3130",x"3332",x"3534",x"3736",x"3938",
--	
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",
--		x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020",x"2020"
--
--	);
--	signal read_addra : std_logic_vector(ADDR_WIDTH-1 downto 0);
--	signal read_addrb : std_logic_vector(ADDR_WIDTH-1 downto 0);
--begin
--	process (ck)
--	begin
--		if (rising_edge(ck)) then
--			if (en = '1') then
--				if (we = '1') then
--					vga_ram(conv_integer(addra)) <= di;
--				end if;
--				read_addra <= addra;
--				read_addrb <= addrb;
--			end if;
--		end if;
--	end process;
--	doa <= vga_ram(conv_integer(read_addra));
--	dob <= vga_ram(conv_integer(read_addrb));
--end Width16;

------------------------------------------------------------------------------------------
--											End of file
--------------------------------------------------------------------------------------------
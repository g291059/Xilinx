----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:33:16 08/05/2008 
-- Design Name: 
-- Module Name:    Rom_t - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE; use IEEE.STD_LOGIC_1164.ALL; use IEEE.STD_LOGIC_ARITH.ALL; use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Rom_t is
	generic ( BUS_WIDTH  : integer range 1 to    8 :=    8;
				 ADDR_WIDTH : integer range 1 to   12 :=   12;
				 ROM_DEPTH	: integer range 1 to 4096 := 3072); 
    Port (  do   : out STD_LOGIC_VECTOR( BUS_WIDTH-1 downto 0);
				addr: in  STD_LOGIC_VECTOR( ADDR_WIDTH-1 downto 0);
            ck	 : in  STD_LOGIC;
				rst : in  STD_LOGIC);
end Rom_t;

architecture Behavioral of Rom_t is

		type romBuff is array (0 to ROM_DEPTH - 1) of std_logic_vector(BUS_WIDTH-1 downto 0);
		constant VGA_ROM : romBuff :=
		(
				x"7E",x"C3",x"99",x"99",x"F3",x"E7",x"E7",x"FF",x"E7",x"E7",x"7E",x"00",	-- x00
				x"00",x"00",x"00",x"76",x"DC",x"00",x"76",x"DC",x"00",x"00",x"00",x"00",
				x"6E",x"D8",x"D8",x"D8",x"D8",x"DE",x"D8",x"D8",x"D8",x"6E",x"00",x"00",
				x"00",x"00",x"00",x"6E",x"DB",x"DB",x"DF",x"D8",x"DB",x"6E",x"00",x"00",
				x"00",x"00",x"10",x"38",x"7C",x"FE",x"7C",x"38",x"10",x"00",x"00",x"00",
				x"88",x"88",x"F8",x"88",x"88",x"00",x"3E",x"08",x"08",x"08",x"08",x"00",
				x"F8",x"80",x"E0",x"80",x"80",x"00",x"3E",x"20",x"38",x"20",x"20",x"00",
				x"78",x"80",x"80",x"80",x"78",x"00",x"3C",x"22",x"3E",x"24",x"22",x"00",
				x"80",x"80",x"80",x"80",x"F8",x"00",x"3E",x"20",x"38",x"20",x"20",x"00",
				x"22",x"88",x"22",x"88",x"22",x"88",x"22",x"88",x"22",x"88",x"22",x"88",
				x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",
				x"EE",x"BB",x"EE",x"BB",x"EE",x"BB",x"EE",x"BB",x"EE",x"BB",x"EE",x"BB",
				x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
				x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
				x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
				x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
				x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",	-- x10
				x"88",x"C8",x"A8",x"98",x"88",x"00",x"20",x"20",x"20",x"20",x"3E",x"00",
				x"88",x"88",x"50",x"50",x"20",x"00",x"3E",x"08",x"08",x"08",x"08",x"00",
				x"00",x"00",x"06",x"0C",x"18",x"30",x"7E",x"00",x"7E",x"00",x"00",x"00",
				x"00",x"00",x"60",x"30",x"18",x"0C",x"7E",x"00",x"7E",x"00",x"00",x"00",
				x"00",x"00",x"06",x"0C",x"FE",x"38",x"FE",x"60",x"C0",x"00",x"00",x"00",
				x"00",x"02",x"0E",x"3E",x"7E",x"FE",x"7E",x"3E",x"0E",x"02",x"00",x"00",
				x"00",x"80",x"E0",x"F0",x"FC",x"FE",x"FC",x"F0",x"E0",x"80",x"00",x"00",
				x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",
				x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"7E",x"3C",x"18",x"00",x"00",
				x"00",x"00",x"00",x"18",x"0C",x"FE",x"0C",x"18",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"30",x"60",x"FE",x"60",x"30",x"00",x"00",x"00",x"00",
				x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"7E",x"3C",x"18",x"00",x"00",
				x"00",x"00",x"00",x"28",x"6C",x"FE",x"6C",x"28",x"00",x"00",x"00",x"00",
				x"00",x"06",x"06",x"36",x"66",x"FE",x"60",x"30",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"C0",x"7C",x"6E",x"6C",x"6C",x"6C",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	-- x20
				x"00",x"18",x"3C",x"3C",x"3C",x"18",x"18",x"00",x"18",x"18",x"00",x"00",
				x"00",x"36",x"36",x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"6C",x"FE",x"6C",x"6C",x"6C",x"FE",x"6C",x"00",x"00",
				x"00",x"10",x"7C",x"D6",x"70",x"38",x"1C",x"D6",x"7C",x"10",x"00",x"00",
				x"00",x"00",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"C6",x"00",x"00",
				x"00",x"38",x"6C",x"38",x"38",x"72",x"FE",x"CC",x"CC",x"76",x"00",x"00",
				x"1C",x"1C",x"0C",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"0C",x"18",x"30",x"30",x"30",x"30",x"30",x"18",x"0C",x"00",x"00",
				x"00",x"30",x"18",x"0C",x"0C",x"0C",x"0C",x"0C",x"18",x"30",x"00",x"00",
				x"00",x"00",x"00",x"6C",x"38",x"FE",x"38",x"6C",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"0C",x"0C",x"18",x"00",
				x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",
				x"00",x"00",x"00",x"06",x"0C",x"18",x"30",x"60",x"C0",x"00",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C6",x"D6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",	-- x30
				x"00",x"18",x"78",x"18",x"18",x"18",x"18",x"18",x"18",x"7E",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"0C",x"18",x"30",x"60",x"C6",x"FE",x"00",x"00",
				x"00",x"7C",x"C6",x"06",x"06",x"3C",x"06",x"06",x"C6",x"7C",x"00",x"00",
				x"00",x"0C",x"1C",x"3C",x"6C",x"CC",x"FE",x"0C",x"0C",x"0C",x"00",x"00",
				x"00",x"FE",x"C0",x"C0",x"C0",x"FC",x"06",x"06",x"C6",x"7C",x"00",x"00",
				x"00",x"7C",x"C6",x"C0",x"C0",x"FC",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"FE",x"C6",x"0C",x"18",x"30",x"30",x"30",x"30",x"30",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C6",x"7C",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C6",x"7E",x"06",x"06",x"C6",x"7C",x"00",x"00",
				x"00",x"00",x"00",x"0C",x"0C",x"00",x"00",x"0C",x"0C",x"00",x"00",x"00",
				x"00",x"00",x"00",x"0C",x"0C",x"00",x"00",x"0C",x"0C",x"0C",x"18",x"00",
				x"00",x"0C",x"18",x"30",x"60",x"C0",x"60",x"30",x"18",x"0C",x"00",x"00",
				x"00",x"00",x"00",x"00",x"FE",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
				x"00",x"60",x"30",x"18",x"0C",x"06",x"0C",x"18",x"30",x"60",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"0C",x"18",x"18",x"00",x"18",x"18",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"DE",x"DE",x"DE",x"DC",x"C0",x"7E",x"00",x"00",
				x"00",x"38",x"6C",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"00",x"00",
				x"00",x"FC",x"66",x"66",x"66",x"7C",x"66",x"66",x"66",x"FC",x"00",x"00",
				x"00",x"3C",x"66",x"C0",x"C0",x"C0",x"C0",x"C0",x"66",x"3C",x"00",x"00",
				x"00",x"F8",x"6C",x"66",x"66",x"66",x"66",x"66",x"6C",x"F8",x"00",x"00",
				x"00",x"FE",x"66",x"60",x"60",x"7C",x"60",x"60",x"66",x"FE",x"00",x"00",
				x"00",x"FE",x"66",x"60",x"60",x"7C",x"60",x"60",x"60",x"F0",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C0",x"C0",x"CE",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"C6",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"C6",x"00",x"00",
				x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"D8",x"D8",x"70",x"00",x"00",
				x"00",x"C6",x"CC",x"D8",x"F0",x"F0",x"D8",x"CC",x"C6",x"C6",x"00",x"00",
				x"00",x"F0",x"60",x"60",x"60",x"60",x"60",x"62",x"66",x"FE",x"00",x"00",
				x"00",x"C6",x"C6",x"EE",x"FE",x"D6",x"D6",x"D6",x"C6",x"C6",x"00",x"00",
				x"00",x"C6",x"C6",x"E6",x"E6",x"F6",x"DE",x"CE",x"CE",x"C6",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"FC",x"66",x"66",x"66",x"7C",x"60",x"60",x"60",x"F0",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"D6",x"7C",x"06",x"00",
				x"00",x"FC",x"66",x"66",x"66",x"7C",x"78",x"6C",x"66",x"E6",x"00",x"00",
				x"00",x"7C",x"C6",x"C0",x"60",x"38",x"0C",x"06",x"C6",x"7C",x"00",x"00",
				x"00",x"7E",x"5A",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"6C",x"38",x"10",x"00",x"00",
				x"00",x"C6",x"C6",x"D6",x"D6",x"D6",x"FE",x"EE",x"C6",x"C6",x"00",x"00",
				x"00",x"C6",x"C6",x"6C",x"38",x"38",x"38",x"6C",x"C6",x"C6",x"00",x"00",
				x"00",x"66",x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"FE",x"C6",x"8C",x"18",x"30",x"60",x"C2",x"C6",x"FE",x"00",x"00",
				x"00",x"7C",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"7C",x"00",x"00",
				x"00",x"00",x"00",x"C0",x"60",x"30",x"18",x"0C",x"06",x"00",x"00",x"00",
				x"00",x"7C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"7C",x"00",x"00",
				x"00",x"18",x"3C",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
				x"1C",x"1C",x"18",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"00",x"E0",x"60",x"60",x"7C",x"66",x"66",x"66",x"66",x"FC",x"00",x"00",
				x"00",x"00",x"00",x"00",x"7C",x"C6",x"C0",x"C0",x"C6",x"7C",x"00",x"00",
				x"00",x"1C",x"0C",x"0C",x"7C",x"CC",x"CC",x"CC",x"CC",x"7E",x"00",x"00",
				x"00",x"00",x"00",x"00",x"7C",x"C6",x"FE",x"C0",x"C6",x"7C",x"00",x"00",
				x"00",x"1C",x"36",x"30",x"30",x"FC",x"30",x"30",x"30",x"78",x"00",x"00",
				x"00",x"00",x"00",x"00",x"76",x"CE",x"C6",x"C6",x"7E",x"06",x"C6",x"7C",
				x"00",x"E0",x"60",x"60",x"6C",x"76",x"66",x"66",x"66",x"E6",x"00",x"00",
				x"00",x"18",x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"00",x"0C",x"0C",x"00",x"1C",x"0C",x"0C",x"0C",x"CC",x"CC",x"78",
				x"00",x"E0",x"60",x"60",x"66",x"6C",x"78",x"6C",x"66",x"E6",x"00",x"00",
				x"00",x"70",x"30",x"30",x"30",x"30",x"30",x"30",x"34",x"18",x"00",x"00",
				x"00",x"00",x"00",x"00",x"6C",x"FE",x"D6",x"D6",x"C6",x"C6",x"00",x"00",
				x"00",x"00",x"00",x"00",x"DC",x"66",x"66",x"66",x"66",x"66",x"00",x"00",
				x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"00",x"00",x"00",x"DC",x"66",x"66",x"66",x"7C",x"60",x"60",x"F0",
				x"00",x"00",x"00",x"00",x"76",x"CC",x"CC",x"CC",x"7C",x"0C",x"0C",x"1E",
				x"00",x"00",x"00",x"00",x"DC",x"66",x"60",x"60",x"60",x"F0",x"00",x"00",
				x"00",x"00",x"00",x"00",x"7C",x"C6",x"70",x"1C",x"C6",x"7C",x"00",x"00",
				x"00",x"30",x"30",x"30",x"FC",x"30",x"30",x"30",x"36",x"1C",x"00",x"00",
				x"00",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",
				x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"6C",x"38",x"10",x"00",x"00",
				x"00",x"00",x"00",x"00",x"C6",x"C6",x"D6",x"D6",x"FE",x"6C",x"00",x"00",
				x"00",x"00",x"00",x"00",x"C6",x"6C",x"38",x"38",x"6C",x"C6",x"00",x"00",
				x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"CE",x"76",x"06",x"C6",x"7C",
				x"00",x"00",x"00",x"00",x"FE",x"8C",x"18",x"30",x"62",x"FE",x"00",x"00",
				x"00",x"0E",x"18",x"18",x"18",x"70",x"18",x"18",x"18",x"0E",x"00",x"00",
				x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",
				x"00",x"70",x"18",x"18",x"18",x"0E",x"18",x"18",x"18",x"70",x"00",x"00",
				x"00",x"76",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"66",x"66",x"00",x"66",x"66",x"66",x"3C",x"18",x"18",x"3C",x"00",x"00",
				x"30",x"18",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",
				x"18",x"30",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",
				x"38",x"6C",x"38",x"00",x"7C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",
				x"76",x"DC",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",
				x"6C",x"6C",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",
				x"38",x"6C",x"38",x"00",x"7C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",
				x"7E",x"D8",x"D8",x"D8",x"D8",x"FE",x"D8",x"D8",x"D8",x"DE",x"00",x"00",
				x"00",x"3C",x"66",x"C0",x"C0",x"C0",x"C6",x"66",x"3C",x"18",x"CC",x"38",
				x"18",x"0C",x"00",x"FE",x"66",x"60",x"7C",x"60",x"66",x"FE",x"00",x"00",
				x"18",x"30",x"00",x"FE",x"66",x"60",x"7C",x"60",x"66",x"FE",x"00",x"00",
				x"38",x"6C",x"00",x"FE",x"66",x"60",x"7C",x"60",x"66",x"FE",x"00",x"00",
				x"6C",x"6C",x"00",x"FE",x"66",x"60",x"7C",x"60",x"66",x"FE",x"00",x"00",
				x"18",x"0C",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"18",x"30",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"3C",x"66",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"66",x"66",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"F8",x"6C",x"66",x"66",x"F6",x"66",x"66",x"6C",x"F8",x"00",x"00",
				x"76",x"DC",x"00",x"C6",x"E6",x"F6",x"DE",x"CE",x"C6",x"C6",x"00",x"00",
				x"30",x"18",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"18",x"30",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"38",x"6C",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"76",x"DC",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"6C",x"6C",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"00",x"00",x"00",x"6C",x"38",x"38",x"6C",x"00",x"00",x"00",x"00",
				x"00",x"7E",x"C6",x"CE",x"DE",x"D6",x"F6",x"E6",x"C6",x"FC",x"00",x"00",
				x"30",x"18",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"18",x"30",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"38",x"6C",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"6C",x"6C",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"0C",x"18",x"00",x"66",x"66",x"66",x"3C",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"F0",x"60",x"7C",x"66",x"66",x"66",x"7C",x"60",x"F0",x"00",x"00",
				x"00",x"7C",x"C6",x"C6",x"C6",x"CC",x"C6",x"C6",x"D6",x"DC",x"80",x"00",
				x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FE",x"00",
				x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"3C",x"3C",x"3C",x"18",
				x"00",x"00",x"10",x"7C",x"D6",x"D0",x"D0",x"D6",x"7C",x"10",x"00",x"00",
				x"00",x"38",x"6C",x"60",x"60",x"F0",x"60",x"66",x"F6",x"6C",x"00",x"00",
				x"00",x"3C",x"62",x"60",x"F8",x"60",x"F8",x"60",x"62",x"3C",x"00",x"00",
				x"00",x"66",x"66",x"3C",x"18",x"7E",x"18",x"3C",x"18",x"18",x"00",x"00",
				x"6C",x"38",x"00",x"7C",x"C6",x"C0",x"7C",x"06",x"C6",x"7C",x"00",x"00",
				x"7C",x"C6",x"C6",x"60",x"7C",x"C6",x"C6",x"7C",x"0C",x"C6",x"C6",x"7C",
				x"00",x"6C",x"38",x"00",x"7C",x"C6",x"70",x"1C",x"C6",x"7C",x"00",x"00",
				x"7E",x"81",x"99",x"A5",x"A1",x"A1",x"A5",x"99",x"81",x"7E",x"00",x"00",
				x"3C",x"6C",x"6C",x"3E",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"36",x"6C",x"D8",x"6C",x"36",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"7E",x"06",x"06",x"06",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",
				x"7E",x"81",x"B9",x"A5",x"A5",x"B9",x"A5",x"A5",x"81",x"7E",x"00",x"00",
				x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"38",x"6C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"7E",x"00",x"00",
				x"00",x"38",x"6C",x"18",x"30",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"38",x"6C",x"18",x"6C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",
				x"6C",x"38",x"00",x"FE",x"C6",x"0C",x"38",x"62",x"C6",x"FE",x"00",x"00",
				x"00",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"F6",x"C0",x"C0",
				x"00",x"7F",x"DB",x"DB",x"DB",x"7B",x"1B",x"1B",x"1B",x"1B",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",
				x"00",x"6C",x"38",x"00",x"FE",x"8C",x"18",x"30",x"62",x"FE",x"00",x"00",
				x"00",x"30",x"70",x"30",x"30",x"78",x"00",x"00",x"00",x"00",x"00",x"00",
				x"38",x"6C",x"6C",x"38",x"00",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"D8",x"6C",x"36",x"6C",x"D8",x"00",x"00",x"00",x"00",
				x"00",x"6E",x"DB",x"DB",x"DF",x"D8",x"D8",x"D9",x"DF",x"6E",x"00",x"00",
				x"00",x"00",x"00",x"00",x"6C",x"DA",x"DE",x"D8",x"DA",x"6C",x"00",x"00",
				x"66",x"66",x"00",x"66",x"66",x"3C",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"00",x"00",x"30",x"30",x"00",x"30",x"30",x"60",x"C6",x"C6",x"7C",
				x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
				x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",
				x"18",x"18",x"18",x"18",x"18",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
				x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
				x"00",x"00",x"00",x"00",x"00",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",
				x"18",x"18",x"18",x"18",x"18",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",
				x"00",x"00",x"00",x"00",x"00",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",
				x"18",x"18",x"18",x"18",x"18",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
				x"18",x"18",x"18",x"18",x"18",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"00",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",
				x"18",x"18",x"18",x"18",x"18",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",
				x"00",x"00",x"00",x"00",x"00",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",
				x"18",x"18",x"18",x"18",x"18",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",
				x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
				x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"7C",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"3F",x"30",x"3F",x"00",x"00",x"00",x"00",x"00",
				x"6C",x"6C",x"6C",x"6C",x"6F",x"60",x"7F",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"7C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"00",x"00",x"00",x"00",x"7F",x"60",x"6F",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"6C",x"6C",x"6C",x"6C",x"6F",x"60",x"6F",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"00",x"00",x"00",x"00",x"FC",x"0C",x"FC",x"00",x"00",x"00",x"00",x"00",
				x"6C",x"6C",x"6C",x"6C",x"EC",x"0C",x"FC",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
				x"6C",x"6C",x"6C",x"6C",x"EF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"FC",x"0C",x"EC",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"6C",x"6C",x"6C",x"6C",x"EC",x"0C",x"EC",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"00",x"00",x"00",x"00",x"FF",x"00",x"EF",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"6C",x"6C",x"6C",x"6C",x"EF",x"00",x"EF",x"6C",x"6C",x"6C",x"6C",x"6C",
				x"60",x"30",x"18",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"18",x"30",x"60",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"30",x"78",x"CC",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"00",x"76",x"DC",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"00",x"6C",x"6C",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"38",x"6C",x"38",x"00",x"78",x"0C",x"7C",x"CC",x"DC",x"76",x"00",x"00",
				x"00",x"00",x"00",x"7E",x"DB",x"1B",x"7F",x"D8",x"DB",x"7E",x"00",x"00",
				x"00",x"00",x"00",x"7C",x"C6",x"C0",x"C0",x"C6",x"7C",x"18",x"6C",x"38",
				x"30",x"18",x"0C",x"00",x"7C",x"C6",x"FE",x"C0",x"C6",x"7C",x"00",x"00",
				x"0C",x"18",x"30",x"00",x"7C",x"C6",x"FE",x"C0",x"C6",x"7C",x"00",x"00",
				x"10",x"38",x"6C",x"00",x"7C",x"C6",x"FE",x"C0",x"C6",x"7C",x"00",x"00",
				x"00",x"6C",x"6C",x"00",x"7C",x"C6",x"FE",x"C0",x"C6",x"7C",x"00",x"00",
				x"60",x"30",x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"0C",x"18",x"30",x"00",x"38",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"18",x"3C",x"66",x"00",x"38",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"00",x"6C",x"6C",x"00",x"38",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",
				x"78",x"30",x"78",x"0C",x"7E",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"76",x"DC",x"00",x"DC",x"66",x"66",x"66",x"66",x"66",x"00",x"00",
				x"60",x"30",x"18",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"0C",x"18",x"30",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"10",x"38",x"6C",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"76",x"DC",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"6C",x"6C",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",
				x"00",x"00",x"18",x"18",x"00",x"7E",x"00",x"18",x"18",x"00",x"00",x"00",
				x"00",x"00",x"00",x"00",x"7E",x"CE",x"DE",x"F6",x"E6",x"FC",x"00",x"00",
				x"C0",x"60",x"30",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",
				x"0C",x"18",x"30",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",
				x"30",x"78",x"CC",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",
				x"00",x"CC",x"CC",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",
				x"0C",x"18",x"30",x"00",x"C6",x"C6",x"C6",x"CE",x"76",x"06",x"C6",x"7C",
				x"00",x"F0",x"60",x"60",x"78",x"6C",x"6C",x"6C",x"78",x"60",x"60",x"F0",
				x"00",x"C6",x"C6",x"00",x"C6",x"C6",x"C6",x"CE",x"76",x"06",x"C6",x"7C"

	);  

begin

	process (ck,rst)
		begin
����� 	if (rst = '1') then
	������	do <= (others => '0');
����� � 	elsif (rising_edge(ck)) then				
				do <= VGA_ROM(conv_integer(addr));
			end if;
		end process;
end Behavioral;

------------------------------------------------------------------------------------------
--		ROM_t2 (16 bit output)
--------------------------------------------------------------------------------------------
library IEEE; use IEEE.STD_LOGIC_1164.ALL; use IEEE.STD_LOGIC_ARITH.ALL; use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Rom_t2 is
	generic ( BUS_WIDTH  : integer range 1 to  16 :=  16;
				 ADDR_WIDTH : integer range 1 to   8 :=   8;
				 ROM_DEPTH	: integer range 1 to 256 := 256); 
    Port (  do   : out STD_LOGIC_VECTOR( BUS_WIDTH-1 downto 0);
				addr: in  STD_LOGIC_VECTOR( ADDR_WIDTH-1 downto 0);
            ck	 : in  STD_LOGIC;
				rst : in  STD_LOGIC);
end Rom_t2;

architecture Behavioral of Rom_t2 is		
	type romBuff is array (0 to ROM_DEPTH - 1) of std_logic_vector(BUS_WIDTH-1 downto 0);
	constant VGA_ROM : romBuff :=
	(
			x"3030",x"3031",x"3032",x"3033",x"3034",x"3035",x"3036",x"3037",	-- 00,01,02,03,04,05,06,07
			x"3038",x"3039",x"3041",x"3042",x"3043",x"3044",x"3045",x"3046",	-- 08,09,0a,0b,0c,0d,0e,0f
			x"3130",x"3131",x"3132",x"3133",x"3134",x"3135",x"3136",x"3137",	-- 10,01,02,03,04,05,06,07
			x"3138",x"3139",x"3141",x"3142",x"3143",x"3144",x"3145",x"3146",	-- 18,09,0a,0b,0c,0d,0e,0f
			x"3230",x"3231",x"3232",x"3233",x"3234",x"3235",x"3236",x"3237",	-- 20,01,02,03,04,05,06,07
			x"3238",x"3239",x"3241",x"3242",x"3243",x"3244",x"3245",x"3246",	-- 28,09,0a,0b,0c,0d,0e,0f
			x"3330",x"3331",x"3332",x"3333",x"3334",x"3335",x"3336",x"3337",	-- 30,01,02,03,04,05,06,07
			x"3338",x"3339",x"3341",x"3342",x"3343",x"3344",x"3345",x"3346",	-- 38,09,0a,0b,0c,0d,0e,0f
			x"3430",x"3431",x"3432",x"3433",x"3434",x"3435",x"3436",x"3437",	-- 40,01,02,03,04,05,06,07
			x"3438",x"3439",x"3441",x"3442",x"3443",x"3444",x"3445",x"3446",	-- 48,09,0a,0b,0c,0d,0e,0f
			x"3530",x"3531",x"3532",x"3533",x"3534",x"3535",x"3536",x"3537",	-- 50,01,02,03,04,05,06,07
			x"3538",x"3539",x"3541",x"3542",x"3543",x"3544",x"3545",x"3546",	-- 58,09,0a,0b,0c,0d,0e,0f
			x"3630",x"3631",x"3632",x"3633",x"3634",x"3635",x"3636",x"3637",	-- 60,01,02,03,04,05,06,07
			x"3638",x"3639",x"3641",x"3642",x"3643",x"3644",x"3645",x"3646",	-- 68,09,0a,0b,0c,0d,0e,0f
			x"3730",x"3731",x"3732",x"3733",x"3734",x"3735",x"3736",x"3737",	-- 70,01,02,03,04,05,06,07
			x"3738",x"3739",x"3741",x"3742",x"3743",x"3744",x"3745",x"3746",	-- 78,09,0a,0b,0c,0d,0e,0f
			x"3830",x"3831",x"3832",x"3833",x"3834",x"3835",x"3836",x"3837",	-- 80,01,02,03,04,05,06,07
			x"3838",x"3839",x"3841",x"3842",x"3843",x"3844",x"3845",x"3846",	-- 88,09,0a,0b,0c,0d,0e,0f
			x"3930",x"3931",x"3932",x"3933",x"3934",x"3935",x"3936",x"3937",	-- 90,01,02,03,04,05,06,07
			x"3938",x"3939",x"3941",x"3942",x"3943",x"3944",x"3945",x"3946",	-- 98,09,0a,0b,0c,0d,0e,0f
			x"4130",x"4131",x"4132",x"4133",x"4134",x"4135",x"4136",x"4137",	-- A0,01,02,03,04,05,06,07
			x"4138",x"4139",x"4141",x"4142",x"4143",x"4144",x"4145",x"4146",	-- A8,09,0a,0b,0c,0d,0e,0f
			x"4230",x"4231",x"4232",x"4233",x"4234",x"4235",x"4236",x"4237",	-- B0,01,02,03,04,05,06,07
			x"4238",x"4239",x"4241",x"4242",x"4243",x"4244",x"4245",x"4246",	-- B8,09,0a,0b,0c,0d,0e,0f
			x"4330",x"4331",x"4332",x"4333",x"4334",x"4335",x"4336",x"4337",	-- C0,01,02,03,04,05,06,07
			x"4338",x"4339",x"4341",x"4342",x"4343",x"4344",x"4345",x"4346",	-- C8,09,0a,0b,0c,0d,0e,0f
			x"4430",x"4431",x"4432",x"4433",x"4434",x"4435",x"4436",x"4437",	-- D0,01,02,03,04,05,06,07
			x"4438",x"4439",x"4441",x"4442",x"4443",x"4444",x"4445",x"4446",	-- D8,09,0a,0b,0c,0d,0e,0f
			x"4530",x"4531",x"4532",x"4533",x"4534",x"4535",x"4536",x"4537",	-- E0,01,02,03,04,05,06,07
			x"4538",x"4539",x"4541",x"4542",x"4543",x"4544",x"4545",x"4546",	-- E8,09,0a,0b,0c,0d,0e,0f
			x"4630",x"4631",x"4632",x"4633",x"4634",x"4635",x"4636",x"4637",	-- F0,01,02,03,04,05,06,07
			x"4638",x"4639",x"4641",x"4642",x"4643",x"4644",x"4645",x"4646"	-- F8,09,0a,0b,0c,0d,0e,0f
	);  

begin

	process (ck,rst)
		begin
����� 	if (rst = '1') then
	������	do <= (others => '0');
����� � 	elsif (rising_edge(ck)) then				
				do <= VGA_ROM(conv_integer(addr));
			end if;
		end process;
end Behavioral;
------------------------------------------------------------------------------------------
--											End of file
--------------------------------------------------------------------------------------------